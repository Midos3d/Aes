module test_bench();

  reg [127:0] in;
  reg [127:0] key;
  reg [127:0] out,fin;
  reg [31:0] R[0:3];
  reg [31:0] t[0:3];
  reg [1:0] bs;
  reg [31:0] rd,rs1,rs2,rdF;
  wire [0:(128*(10+1))-1 ] fullkeys;
  int i;
keyExpansion  ke (key,fullkeys);
  aes32esmi aes (bs,rs1,rs2,rd);
  aes32esi aesF (bs,rs1,rs2,rdF);
  initial 
    begin
      key =128'h_000102030405060708090a0b0c0d0e0f;
      in = 128'h_00112233445566778899aabbccddeeff;
      #1
      out = key^in;
      #1
      t[0]=out[127:96];
      t[1]=out[95:64];
      t[2]=out[63:32];
      t[3]=out[31:0];
      
      for(i=1;i<10;i++)
        begin
          #1
          R[0]=fullkeys[128*i +:32];
          R[1]=fullkeys[(128*i+32) +:32];
          R[2]=fullkeys[(128*i+64)+:32];
          R[3]=fullkeys[(128*i+96)+:32];
    
      #1
      /////////////////row 1
          bs=0;
      rs2=t[0];
      rs1=R[0];
      #1
      R[0]=rd;
      #1
          bs=1;
      rs2=t[1];
      rs1=R[0];
      #1
      R[0]=rd;
      #1
          bs=2;
      rs2=t[2];
      rs1=R[0];
      #1
      R[0]=rd;
      #1
          bs=3;
      rs2=t[3];
      rs1=R[0];
      #1
      R[0]=rd;
      #1
      
      
       /////////////////row 2
      
      bs=0;
      rs2=t[1];
      rs1=R[1];
      #1
      R[1]=rd;
      #1
          bs=1;
      rs2=t[2];
      rs1=R[1];
      #1
      R[1]=rd;
      #1
          bs=2;
      rs2=t[3];
      rs1=R[1];
      #1
      R[1]=rd;
      #1
          bs=3;
      rs2=t[0];
      rs1=R[1];
      #1
      R[1]=rd;
      #1
      
       /////////////////row 3
      
           bs=0;
      rs2=t[2];
      rs1=R[2];
      #1
      R[2]=rd;
      #1
          bs=1;
      rs2=t[3];
      rs1=R[2];
      #1
      R[2]=rd;
      #1
          bs=2;
      rs2=t[0];
      rs1=R[2];
      #1
      R[2]=rd;
      #1
          bs=3;
      rs2=t[1];
      rs1=R[2];
      #1
      R[2]=rd;
      #1
      
      
      
       /////////////////row 4
      
            bs=0;
      rs2=t[3];
      rs1=R[3];
      #1
      R[3]=rd;
      #1
          bs=1;
      rs2=t[0];
      rs1=R[3];
      #1
      R[3]=rd;
      #1
          bs=2;
      rs2=t[1];
      rs1=R[3];
      #1
      R[3]=rd;
      #1
          bs=3;
      rs2=t[2];
      rs1=R[3];
      #1
      R[3]=rd;
     #1
          t[0]=R[0];
          t[1]=R[1];
          t[2]=R[2];
          t[3]=R[3];

        end
       #1
      R[0]=fullkeys[128*10 +:32];
      R[1]=fullkeys[(128*10+32) +:32];
      R[2]=fullkeys[(128*10+64)+:32];
      R[3]=fullkeys[(128*10+96)+:32];
      
      
       #1
      /////////////////row 1
          bs=0;
      rs2=t[0];
      rs1=R[0];
      #1
      R[0]=rdF;
      #1
          bs=1;
      rs2=t[1];
      rs1=R[0];
      #1
      R[0]=rdF;
      #1
          bs=2;
      rs2=t[2];
      rs1=R[0];
      #1
      R[0]=rdF;
      #1
          bs=3;
      rs2=t[3];
      rs1=R[0];
      #1
      R[0]=rdF;
      #1
      
      
       /////////////////row 2
      
      bs=0;
      rs2=t[1];
      rs1=R[1];
      #1
      R[1]=rdF;
      #1
          bs=1;
      rs2=t[2];
      rs1=R[1];
      #1
      R[1]=rdF;
      #1
          bs=2;
      rs2=t[3];
      rs1=R[1];
      #1
      R[1]=rdF;
      #1
          bs=3;
      rs2=t[0];
      rs1=R[1];
      #1
      R[1]=rdF;
      #1
      
       /////////////////row 3
      
           bs=0;
      rs2=t[2];
      rs1=R[2];
      #1
      R[2]=rdF;
      #1
          bs=1;
      rs2=t[3];
      rs1=R[2];
      #1
      R[2]=rdF;
      #1
          bs=2;
      rs2=t[0];
      rs1=R[2];
      #1
      R[2]=rdF;
      #1
          bs=3;
      rs2=t[1];
      rs1=R[2];
      #1
      R[2]=rdF;
      #1
      
      
      
       /////////////////row 4
      
            bs=0;
      rs2=t[3];
      rs1=R[3];
      #1
      R[3]=rdF;
      #1
          bs=1;
      rs2=t[0];
      rs1=R[3];
      #1
      R[3]=rdF;
      #1
          bs=2;
      rs2=t[1];
      rs1=R[3];
      #1
      R[3]=rdF;
      #1
          bs=3;
      rs2=t[2];
      rs1=R[3];
      #1
      R[3]=rdF;
     #1
      
       fin ={R[0],R[1],R[2],R[3]};
      #1
      $display("%0h", fin);
      
    end

  
  
  
  

  
endmodule